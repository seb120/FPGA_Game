//-------------------------------------------------------------------------
//      lab7_usb.sv                                                      --
//      Christine Chen                                                   --
//      Fall 2014                                                        --
//                                                                       --
//      Fall 2014 Distribution                                           --
//                                                                       --
//      For use with ECE 385 Lab 7                                       --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------


module  lab7_usb 		( input         Clk,
                                     Reset,
							  output [6:0]  HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7,
							  output [8:0]  LEDG,
							  output [17:0] LEDR,
							  // VGA Interface 
                       output [7:0]  Red,
							                Green,
												 Blue,
							  output        VGA_clk,
							                sync,
												 blank,
												 vs,
												 hs,
							  // CY7C67200 Interface
							  inout [15:0]  OTG_DATA,						//	CY7C67200 Data bus 16 Bits
							  output [1:0]  OTG_ADDR,						//	CY7C67200 Address 2 Bits
							  output        OTG_CS_N,						//	CY7C67200 Chip Select
												 OTG_RD_N,						//	CY7C67200 Write
												 OTG_WR_N,						//	CY7C67200 Read
												 OTG_RST_N,						//	CY7C67200 Reset
							  input			 OTG_INT,						//	CY7C67200 Interrupt
							  // SDRAM Interface for Nios II Software
							  output [12:0] sdram_wire_addr,				// SDRAM Address 13 Bits
							  inout [31:0]  sdram_wire_dq,				// SDRAM Data 32 Bits
							  output [1:0]  sdram_wire_ba,				// SDRAM Bank Address 2 Bits
							  output [3:0]  sdram_wire_dqm,				// SDRAM Data Mast 4 Bits
							  output			 sdram_wire_ras_n,			// SDRAM Row Address Strobe
							  output			 sdram_wire_cas_n,			// SDRAM Column Address Strobe
							  output			 sdram_wire_cke,				// SDRAM Clock Enable
							  output			 sdram_wire_we_n,				// SDRAM Write Enable
							  output			 sdram_wire_cs_n,				// SDRAM Chip Select
							  output			 sdram_clk						// SDRAM Clock
											);
    
    logic Reset_h, vssig;
	 logic [2:0]pacstatesig;
    logic [9:0] drawxsig, drawysig, pacmanxsig, pacmanysig, spritesizesig, blue_ghostxsig, blue_ghostysig, chXsig, chYsig, oneXsig, oneYsig, twoXsig, twoYsig;
	 logic [9:0] s1Xsig, s1Ysig, c1Xsig, c1Ysig, o1Xsig, o1Ysig, r1Xsig, r1Ysig, e1Xsig, e1Ysig, lvlsig;
	 logic [7:0] keycode;
	 logic reset1, chOnsig, ressig;
	 logic [7:0] scoreval;
    assign {Reset_h}=~ (Reset);  // The push buttons are active low
	 assign OTG_FSPEED = 1'bz;
	 assign OTG_LSPEED = 1'bz;
	    
	 usb_system usbsys_instance(
										 .clk_clk(Clk),         
										 .reset_reset_n(1'b1),   
										 .sdram_wire_addr(sdram_wire_addr), 
										 .sdram_wire_ba(sdram_wire_ba),   
										 .sdram_wire_cas_n(sdram_wire_cas_n),
										 .sdram_wire_cke(sdram_wire_cke),  
										 .sdram_wire_cs_n(sdram_wire_cs_n), 
										 .sdram_wire_dq(sdram_wire_dq),   
										 .sdram_wire_dqm(sdram_wire_dqm),  
										 .sdram_wire_ras_n(sdram_wire_ras_n),
										 .sdram_wire_we_n(sdram_wire_we_n), 
										 .sdram_out_clk_clk(sdram_clk),
										 .keycode_export(keycode),  
										 .usb_DATA(OTG_DATA),    
										 .usb_ADDR(OTG_ADDR),    
										 .usb_RD_N(OTG_RD_N),    
										 .usb_WR_N(OTG_WR_N),    
										 .usb_CS_N(OTG_CS_N),    
										 .usb_RST_N(OTG_RST_N),   
										 .usb_INT(OTG_INT) );
	
    vga_controller vgasync_instance(.*,
	                                 .Clk(Clk),
											   .Reset(Reset_h),
											   .pixel_clk(VGA_clk),
											   .DrawX(drawxsig),
								 			   .DrawY(drawysig) );
   
    Game_entity_table pm_instance(.Reset(Reset_h),
	                    .frame_clk(vs),    // Vertical Sync used as an "ad hoc" 60 Hz clock signal
	                    .key(keycode),
							  .pacmanX(pacmanxsig),  // (This is why we registered it in the vga controller!)
							  .pacmanY(pacmanysig),
							  .pacmanState(pacstatesig),
							  .blue_ghostX(blue_ghostxsig),
							  .blue_ghostY(blue_ghostysig),
							  .ch_X(chXsig),
							  .ch_Y(chYsig),
							  .ch_on(chOnsig),
							  .res(ressig),
							  .onescoreX(oneXsig), 
							  .onescoreY(oneYsig),
							  .twoscoreX(twoXsig),
							  .twoscoreY(twoYsig),
							  .s1X(s1Xsig), 
							  .s1Y(s1Ysig), 
							  .c1X(c1Xsig), 
							  .c1Y(c1Ysig), 
							  .o1X(o1Xsig), 
							  .o1Y(o1Ysig), 
							  .r1X(r1Xsig), 
							  .r1Y(r1Ysig), 
							  .e1X(e1Xsig), 
							  .e1Y(e1Ysig),
							  .lvl(lvlsig),
							  .score(scoreval),
							  .Size(spritesizesig));
							  
   
    color_mapper color_instance(.*,
	                             .pacmanX(pacmanxsig),
		 								  .pacmanY(pacmanysig),
										  .pacState(pacstatesig),
										  .blue_ghostX(blue_ghostxsig),
		 								  .blue_ghostY(blue_ghostysig),
		 								  .DrawX(drawxsig),
		 								  .DrawY(drawysig),
										  .ch_X(chXsig),
										  .ch_Y(chYsig),
							           .ch_on(chOnsig),
										  .onescoreX(oneXsig),
										  .onescoreY(oneYsig),
										  .twoscoreX(twoXsig),
										  .twoscoreY(twoYsig),
										  .s1X(s1Xsig), 
										  .s1Y(s1Ysig), 
										  .c1X(c1Xsig), 
										  .c1Y(c1Ysig), 
										  .o1X(o1Xsig), 
										  .o1Y(o1Ysig), 
										  .r1X(r1Xsig), 
										  .r1Y(r1Ysig), 
										  .e1X(e1Xsig), 
										  .e1Y(e1Ysig),
										  .lvl(lvlsig),
										  .res(ressig),
										  .score(scoreval),
										  .sprite_size(spritesizesig) );
	 

	 HexDriver hex_inst_0 (keycode[3:0], HEX0);
	 HexDriver hex_inst_1 (keycode[7:4], HEX1);
    

	 /**************************************************************************************
	    ATTENTION! Please answer the following quesiton in your lab report! Points will be allocated for the answers!
		 Hidden Question #1/2:
          What are the advantages and/or disadvantages of using a USB interface over PS/2 interface to
			 connect to the keyboard? List any two.  Give an answer in your Post-Lab.
     **************************************************************************************/
endmodule
