library verilog;
use verilog.vl_types.all;
entity altera_avalon_dc_fifo is
    generic(
        SYMBOLS_PER_BEAT: integer := 1;
        BITS_PER_SYMBOL : integer := 8;
        FIFO_DEPTH      : integer := 16;
        CHANNEL_WIDTH   : integer := 0;
        ERROR_WIDTH     : integer := 0;
        USE_PACKETS     : integer := 0;
        USE_IN_FILL_LEVEL: integer := 0;
        USE_OUT_FILL_LEVEL: integer := 0;
        WR_SYNC_DEPTH   : integer := 2;
        RD_SYNC_DEPTH   : integer := 2;
        STREAM_ALMOST_FULL: integer := 0;
        STREAM_ALMOST_EMPTY: integer := 0;
        BACKPRESSURE_DURING_RESET: integer := 0;
        LOOKAHEAD_POINTERS: integer := 0;
        PIPELINE_POINTERS: integer := 0;
        USE_SPACE_AVAIL_IF: integer := 0
    );
    port(
        in_clk          : in     vl_logic;
        in_reset_n      : in     vl_logic;
        out_clk         : in     vl_logic;
        out_reset_n     : in     vl_logic;
        in_data         : in     vl_logic_vector;
        in_valid        : in     vl_logic;
        in_ready        : out    vl_logic;
        in_startofpacket: in     vl_logic;
        in_endofpacket  : in     vl_logic;
        in_empty        : in     vl_logic_vector;
        in_error        : in     vl_logic_vector;
        in_channel      : in     vl_logic_vector;
        out_data        : out    vl_logic_vector;
        out_valid       : out    vl_logic;
        out_ready       : in     vl_logic;
        out_startofpacket: out    vl_logic;
        out_endofpacket : out    vl_logic;
        out_empty       : out    vl_logic_vector;
        out_error       : out    vl_logic_vector;
        out_channel     : out    vl_logic_vector;
        in_csr_address  : in     vl_logic;
        in_csr_write    : in     vl_logic;
        in_csr_read     : in     vl_logic;
        in_csr_readdata : out    vl_logic_vector(31 downto 0);
        in_csr_writedata: in     vl_logic_vector(31 downto 0);
        out_csr_address : in     vl_logic;
        out_csr_write   : in     vl_logic;
        out_csr_read    : in     vl_logic;
        out_csr_readdata: out    vl_logic_vector(31 downto 0);
        out_csr_writedata: in     vl_logic_vector(31 downto 0);
        almost_full_valid: out    vl_logic;
        almost_full_data: out    vl_logic;
        almost_empty_valid: out    vl_logic;
        almost_empty_data: out    vl_logic;
        space_avail_data: out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of SYMBOLS_PER_BEAT : constant is 1;
    attribute mti_svvh_generic_type of BITS_PER_SYMBOL : constant is 1;
    attribute mti_svvh_generic_type of FIFO_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of CHANNEL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ERROR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of USE_PACKETS : constant is 1;
    attribute mti_svvh_generic_type of USE_IN_FILL_LEVEL : constant is 1;
    attribute mti_svvh_generic_type of USE_OUT_FILL_LEVEL : constant is 1;
    attribute mti_svvh_generic_type of WR_SYNC_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of RD_SYNC_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of STREAM_ALMOST_FULL : constant is 1;
    attribute mti_svvh_generic_type of STREAM_ALMOST_EMPTY : constant is 1;
    attribute mti_svvh_generic_type of BACKPRESSURE_DURING_RESET : constant is 1;
    attribute mti_svvh_generic_type of LOOKAHEAD_POINTERS : constant is 1;
    attribute mti_svvh_generic_type of PIPELINE_POINTERS : constant is 1;
    attribute mti_svvh_generic_type of USE_SPACE_AVAIL_IF : constant is 1;
end altera_avalon_dc_fifo;
