module sprite_table ( input [9:0]	addr,
							 output [63:0]	data
					 );
			
	parameter ADDR_WIDTH = 10;
	parameter DATA_WIDTH =  64;
	logic [ADDR_WIDTH-1:0] addr_reg;
	
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
			//code 0000000000 blk box
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 2
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 3
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 4
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 5
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 6
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 7
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 8
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 9
        64'b0000000000000000000000000000000000000000000000000000000000000000, // a
        64'b0000000000000000000000000000000000000000000000000000000000000000, // b
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  // code 0000000000 pig
		  64'b0000000000000001000100000000000000000000000000010001000000000000, // 0
        64'b0000000000000001001000100001000100010001001000100001000000000000, // 1
        64'b0000000000000000000100100010001000100010001000010000000000000000, // 2
        64'b0000000000000000000100100010001000100010001000010000000000000000, // 3
        64'b0000000000000000000000010010001000100010000100000000000000000000, // 4
        64'b0000000000000000000100010010001000100010000100010000000000000000, // 5
        64'b0000000000000001001000100010001000100010001000100001000000000000, // 6
        64'b0000000000000001001000100010001000100010001000100001000000000000, // 7
        64'b0000000000000001001000100010001000100010001000100001000000000000, // 8
        64'b0000000000000001001000100010011001100001001000100001000000000000, // 9
        64'b0000000000000001001000100010000101010001001000100001000000000000, // a
        64'b0000000000000000000100100010000101100110001000010000000000000000, // b
        64'b0000000000000000000100100010001000100010001000010000000000000000, // c
        64'b0000000000000000000100010001000100010001000100010000000000000000, // d
        64'b0000000000000000000000100000000000000000001000000000000000000000, // e
        64'b0000000000000000000001000000000000000000010000000000000000000000, // f
         // code 0000010000 chicken
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  // code 0000100000 shit
		  64'b0000000000000000000000000000101100000000000000000000000000000000, // 0
        64'b0000000000000000000000001011110010110000000000000000000000000000, // 1
        64'b0000000000000000000010111110110011001011000000000000000000000000, // 2
        64'b0000000000000000101111101101110111001100101100000000000000000000, // 3
        64'b0000000000000000101110111101110111011011101100000000000000000000, // 4
        64'b0000000010111011111011101101110111011100110010111011000000000000, // 5
        64'b0000101111101110110111011101110111011101110111001100101100000000, // 6
        64'b1011101110111101110111011101110011011101110111001011101110110000, // 7
        64'b1011111011101101110111011101111011001100110010111100110011001011, // 8
        64'b1011111011011110111011011101110111101110110111011100110011001011, // 9
        64'b1011111011011101110111101110110111011101110111011101110011001011, // a
        64'b1011111011011101110111011101110011011101110111011101110010111011, // b
        64'b0000101111001101110111011101111011001100110011001100101110110000, // c
        64'b0000101110111100110011011101110111101110110111011011101100000000, // d
        64'b0000000000001011101110111011101110111011101110110000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  // code 0000110000 cow
		  64'b0000000010111011000000001011000000000000000000000000000000000000, // 0
        64'b0000101101110111101110110111101100001011101110111011000000000000, // 1
        64'b0000101101110111011111011011101110111101110111010111101110110000, // 2
        64'b0000000010110111011101110111101111011101110111010111101100001011, // 3
        64'b0000000010110111101101111011011101111101110101111101101110110000, // 4
        64'b0000000010110111101101111011011101111101110101111101110110110000, // 5
        64'b0000101101110111011101110111011101111101110101110111011110110000, // 6
        64'b1011011101110111011101110111011111011101110111010111011110110000, // 7
        64'b1011011101110111011101110111110111011101110111011101011110110000, // 8
        64'b1011111111111111111110110111110101111101011111010111011110110000, // 9
        64'b0000101110111111101101110111011101110111011101110111101100000000, // a
        64'b0000000010111011011101110111101101110111101101111011000000000000, // b
        64'b0000000010111011101101110111101110111011000010111011000000000000, // c
        64'b0000000010111011000010111011101100000000000010111011000000000000, // d
        64'b0000000000000000000000001011101100000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  // code 0001000000 sheep
		  64'b0000000000000000000000000000000000000000000000000000000000000000, // 0
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1
        64'b0000000000000000000010111011101110110000101110111011101100000000, // 2
        64'b0000000000000000101101110111011110111011101101110111101110110000, // 3
        64'b0000000010111011101101110111011101110111011101110111011110111011, // 4
        64'b0000101110111011101101110111101101110111011101110111011101111011, // 5
        64'b1011101101111011101110110111011110110111101101110111011101111011, // 6
        64'b1011101110111011011110110111011110110111011110110111011110111011, // 7
        64'b1011101110110111011101110111101101110111011110110111011110110000, // 8
        64'b0000101110111011101101110111011101110111011110110111011110111011, // 9
        64'b0000000000000000101101110111011101110111101101110111011101111011, // a
        64'b0000000000000000101101110111011101110111011101110111011101111011, // b
        64'b0000000000000000101110110111011110111011011101111011011110110000, // c
        64'b0000000000000000000010111011101100000000101110110000101100000000, // d
        64'b0000000000000000000010110000101100000000000010110000101100000000, // e
        64'b0000000000000000000010110000101100000000000010110000101100000000, // f
		  // code 0001010000 '0'
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1
        64'b0000111111111111111111110000000000000000000000000000000000000000, // 2  *****
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 3 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 4 **   **
        64'b1111111100000000111111111111000000000000000000000000000000000000, // 5 **  ***
        64'b1111111100001111111111111111000000000000000000000000000000000000, // 6 ** ****
        64'b1111111111111111000011111111000000000000000000000000000000000000, // 7 **** **
        64'b1111111111110000000011111111000000000000000000000000000000000000, // 8 ***  **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 9 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // a **   **
        64'b0000111111111111111111110000000000000000000000000000000000000000, // b  *****
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  // code 0001100000 '1'
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 2
        64'b0000000011111111111100000000000000000000000000000000000000000000, // 3
        64'b0000111111111111111100000000000000000000000000000000000000000000, // 4    **
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 5   ***
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 6  ****
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 7    **
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 8    **
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 9    **
        64'b0000000000001111111100000000000000000000000000000000000000000000, // a    **
        64'b0000111111111111111111111111000000000000000000000000000000000000, // b    **
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c    **
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d  ******
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
		  		  // code 0001110000 '2'
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b0000111111111111111111110000000000000000000000000000000000000000, // 2  *****
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 3 **   **
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 4      **
        64'b0000000000000000111111110000000000000000000000000000000000000000, // 5     **
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 6    **
        64'b0000000011111111000000000000000000000000000000000000000000000000, // 7   **
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 8  **
        64'b1111111100000000000000000000000000000000000000000000000000000000, // 9 **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // a **   **
        64'b1111111111111111111111111111000000000000000000000000000000000000, // b *******
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0010000000 3
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b0000111111111111111111110000000000000000000000000000000000000000, // 2  *****
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 3 **   **
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 4      **
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 5      **
        64'b0000000011111111111111110000000000000000000000000000000000000000, // 6   ****
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 7      **
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 8      **
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 9      **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // a **   **
        64'b0000111111111111111111110000000000000000000000000000000000000000, // b  *****
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  // code 0010010000 4
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b0000000000000000111111110000000000000000000000000000000000000000, // 2     **
        64'b0000000000001111111111110000000000000000000000000000000000000000, // 3    ***
        64'b0000000011111111111111110000000000000000000000000000000000000000, // 4   ****
        64'b0000111111110000111111110000000000000000000000000000000000000000, // 5  ** **
        64'b1111111100000000111111110000000000000000000000000000000000000000, // 6 **  **
        64'b1111111111111111111111111111000000000000000000000000000000000000, // 7 *******
        64'b0000000000000000111111110000000000000000000000000000000000000000, // 8     **
        64'b0000000000000000111111110000000000000000000000000000000000000000, // 9     **
        64'b0000000000000000111111110000000000000000000000000000000000000000, // a     **
        64'b0000000000001111111111111111000000000000000000000000000000000000, // b    ****
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  // code 0010100000 5
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b1111111111111111111111111111000000000000000000000000000000000000, // 2 *******
        64'b1111111100000000000000000000000000000000000000000000000000000000, // 3 **
        64'b1111111100000000000000000000000000000000000000000000000000000000, // 4 **
        64'b1111111100000000000000000000000000000000000000000000000000000000, // 5 **
        64'b1111111111111111111111110000000000000000000000000000000000000000, // 6 ******
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 7      **
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 8      **
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 9      **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // a **   **
        64'b0000111111111111111111110000000000000000000000000000000000000000, // b  *****
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0010110000 6
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b0000000011111111111100000000000000000000000000000000000000000000, // 2   ***
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 3  **
        64'b1111111100000000000000000000000000000000000000000000000000000000, // 4 **
        64'b1111111100000000000000000000000000000000000000000000000000000000, // 5 **
        64'b1111111111111111111111110000000000000000000000000000000000000000, // 6 ******
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 7 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 8 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 9 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // a **   **
        64'b0000111111111111111111110000000000000000000000000000000000000000, // b  *****
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0011000000 7
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b1111111111111111111111111111000000000000000000000000000000000000, // 2 *******
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 3 **   **
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 4      **
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 5      **
        64'b0000000000000000111111110000000000000000000000000000000000000000, // 6     **
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 7    **
        64'b0000000011111111000000000000000000000000000000000000000000000000, // 8   **
        64'b0000000011111111000000000000000000000000000000000000000000000000, // 9   **
        64'b0000000011111111000000000000000000000000000000000000000000000000, // a   **
        64'b0000000011111111000000000000000000000000000000000000000000000000, // b   **
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0011010000 8
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b0000111111111111111111110000000000000000000000000000000000000000, // 2  *****
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 3 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 4 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 5 **   **
        64'b0000111111111111111111110000000000000000000000000000000000000000, // 6  *****
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 7 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 8 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 9 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // a **   **
        64'b0000111111111111111111110000000000000000000000000000000000000000, // b  *****
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0011100000 9
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b0000111111111111111111000000000000000000000000000000000000000000, // 2  *****
        64'b1111111100000000001111111100000000000000000000000000000000000000, // 3 **   **
        64'b1111111100000000001111111100000000000000000000000000000000000000, // 4 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 5 **   **
        64'b0000111111111111111111111111000000000000000000000000000000000000, // 6  ******
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 7      **
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 8      **
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 9      **
        64'b0000000000000000111111110000000000000000000000000000000000000000, // a     **
        64'b0000111111111111111100000000000000000000000000000000000000000000, // b  ****
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0011110000 A
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b0000000000001111000000000000000000000000000000000000000000000000, // 2    *
        64'b0000000011111111111100000000000000000000000000000000000000000000, // 3   ***
        64'b0000111111110000111111110000000000000000000000000000000000000000, // 4  ** **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 5 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 6 **   **
        64'b1111111111111111111111111111000000000000000000000000000000000000, // 7 *******
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 8 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 9 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // a **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // b **   **
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0100000000 C
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b0000000011111111111111110000000000000000000000000000000000000000, // 2   ****
        64'b0000111111110000000011111111000000000000000000000000000000000000, // 3  **  **
        64'b1111111100000000000000001111000000000000000000000000000000000000, // 4 **    *
        64'b1111111100000000000000000000000000000000000000000000000000000000, // 5 **
        64'b1111111100000000000000000000000000000000000000000000000000000000, // 6 **
        64'b1111111100000000000000000000000000000000000000000000000000000000, // 7 **
        64'b1111111100000000000000000000000000000000000000000000000000000000, // 8 **
        64'b1111111100000000000000001111000000000000000000000000000000000000, // 9 **    *
        64'b0000111111110000000011111111000000000000000000000000000000000000, // a  **  **
        64'b0000000011111111111111110000000000000000000000000000000000000000, // b   ****
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0100010000 E
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b1111111111111111111111111111000000000000000000000000000000000000, // 2 *******
        64'b0000111111110000000011111111000000000000000000000000000000000000, // 3  **  **
        64'b0000111111110000000000001111000000000000000000000000000000000000, // 4  **   *
        64'b0000111111110000111100000000000000000000000000000000000000000000, // 5  ** *
        64'b0000111111111111111100000000000000000000000000000000000000000000, // 6  ****
        64'b0000111111110000111100000000000000000000000000000000000000000000, // 7  ** *
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 8  **
        64'b0000111111110000000000001111000000000000000000000000000000000000, // 9  **   *
        64'b0000111111110000000011111111000000000000000000000000000000000000, // a  **  **
        64'b1111111111111111111111111111000000000000000000000000000000000000, // b *******
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0100100000 G
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b0000000011111111111111110000000000000000000000000000000000000000, // 2   ****
        64'b0000111111110000000011111111000000000000000000000000000000000000, // 3  **  **
        64'b1111111100000000000000001111000000000000000000000000000000000000, // 4 **    *
        64'b1111111100000000000000000000000000000000000000000000000000000000, // 5 **
        64'b1111111100000000000000000000000000000000000000000000000000000000, // 6 **
        64'b1111111100001111111111111111000000000000000000000000000000000000, // 7 ** ****
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 8 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 9 **   **
        64'b0000111111110000000011111111000000000000000000000000000000000000, // a  **  **
        64'b0000000011111111111100001111000000000000000000000000000000000000, // b   *** *
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0100110000 M
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b1111111100000000000000001111111100000000000000000000000000000000, // 2 **    **
        64'b1111111111110000000011111111111100000000000000000000000000000000, // 3 ***  ***
        64'b1111111111111111111111111111111100000000000000000000000000000000, // 4 ********
        64'b1111111111111111111111111111111100000000000000000000000000000000, // 5 ********
        64'b1111111100001111111100001111111100000000000000000000000000000000, // 6 ** ** **
        64'b1111111100000000000000001111111100000000000000000000000000000000, // 7 **    **
        64'b1111111100000000000000001111111100000000000000000000000000000000, // 8 **    **
        64'b1111111100000000000000001111111100000000000000000000000000000000, // 9 **    **
        64'b1111111100000000000000001111111100000000000000000000000000000000, // a **    **
        64'b1111111100000000000000001111111100000000000000000000000000000000, // b **    **
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0101000000 N
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 2 **   **
        64'b1111111111110000000011111111000000000000000000000000000000000000, // 3 ***  **
        64'b1111111111111111000011111111000000000000000000000000000000000000, // 4 **** **
        64'b1111111111111111111111111111000000000000000000000000000000000000, // 5 *******
        64'b1111111100001111111111111111000000000000000000000000000000000000, // 6 ** ****
        64'b1111111100000000111111111111000000000000000000000000000000000000, // 7 **  ***
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 8 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 9 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // a **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // b **   **
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0101010000 O
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b0000111111111111111111110000000000000000000000000000000000000000, // 2  *****
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 3 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 4 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 5 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 6 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 7 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 8 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 9 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // a **   **
        64'b0000111111111111111111110000000000000000000000000000000000000000, // b  *****
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0101100000 R
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b1111111111111111111111110000000000000000000000000000000000000000, // 2 ******
        64'b0000111111110000000011111111000000000000000000000000000000000000, // 3  **  **
        64'b0000111111110000000011111111000000000000000000000000000000000000, // 4  **  **
        64'b0000111111110000000011111111000000000000000000000000000000000000, // 5  **  **
        64'b0000111111111111111111110000000000000000000000000000000000000000, // 6  *****
        64'b0000111111110000111111110000000000000000000000000000000000000000, // 7  ** **
        64'b0000111111110000000011111111000000000000000000000000000000000000, // 8  **  **
        64'b0000111111110000000011111111000000000000000000000000000000000000, // 9  **  **
        64'b0000111111110000000011111111000000000000000000000000000000000000, // a  **  **
        64'b1111111111110000000011111111000000000000000000000000000000000000, // b ***  **
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0101110000 S
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b0000111111111111111111110000000000000000000000000000000000000000, // 2  *****
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 3 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 4 **   **
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 5  **
        64'b0000000011111111111100000000000000000000000000000000000000000000, // 6   ***
        64'b0000000000000000111111110000000000000000000000000000000000000000, // 7     **
        64'b0000000000000000000011111111000000000000000000000000000000000000, // 8      **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // 9 **   **
        64'b1111111100000000000011111111000000000000000000000000000000000000, // a **   **
        64'b0000111111111111111111110000000000000000000000000000000000000000, // b  *****
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0110000000 T
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b1111111111111111111111111111111100000000000000000000000000000000, // 2 ********
        64'b1111111100001111111100001111111100000000000000000000000000000000, // 3 ** ** **
        64'b1111000000001111111100000000111100000000000000000000000000000000, // 4 *  **  *
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 5    **
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 6    **
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 7    **
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 8    **
        64'b0000000000001111111100000000000000000000000000000000000000000000, // 9    **
        64'b0000000000001111111100000000000000000000000000000000000000000000, // a    **
        64'b0000000011111111111111110000000000000000000000000000000000000000, // b   ****
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0110010000 V
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b1111111100000000000000001111111100000000000000000000000000000000, // 2 **    **
        64'b1111111100000000000000001111111100000000000000000000000000000000, // 3 **    **
        64'b1111111100000000000000001111111100000000000000000000000000000000, // 4 **    **
        64'b1111111100000000000000001111111100000000000000000000000000000000, // 5 **    **
        64'b1111111100000000000000001111111100000000000000000000000000000000, // 6 **    **
        64'b1111111100000000000000001111111100000000000000000000000000000000, // 7 **    **
        64'b1111111100000000000000001111111100000000000000000000000000000000, // 8 **    **
        64'b0000111111110000000011111111000000000000000000000000000000000000, // 9  **  **
        64'b0000000011111111111111110000000000000000000000000000000000000000, // a   ****
        64'b0000000000001111111100000000000000000000000000000000000000000000, // b    **
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0110100000 tree
		  64'b0000000000000000000010111011101100001011101110110000000000000000, // 0
        64'b0000000000001011101110110000101110111011000010111011000000000000, // 1
        64'b0000000000001011000000000000000000000000000000001011101100000000, // 2
        64'b0000000010111011000011000000000000000000000011000000101100000000, // 3
        64'b0000000010110000110000000000000000000000000011000000101100000000, // 4
        64'b0000000010110000000000000000000000000000000011000000101100000000, // 5
        64'b0000000010111011000000000000000000000000110000001011101100000000, // 6
        64'b0000000000001011101100000000000000000000000010111011000000000000, // 7
        64'b0000000000000000101110111011101110111011101110110000000000000000, // 8
        64'b0000000000000000000000001101111011101100000000000000000000000000, // 9
        64'b0000000000000000000000001101111011001100000000000000000000000000, // a
        64'b0000000000000000000000001101111011001101000000000000000000000000, // b
        64'b0000000000000000000011011110111011001110110100000000000000000000, // c
        64'b0000000000000000000011011110110011001101110100000000000000000000, // d
        64'b0000000000000000000011011100110011101101110100000000000000000000, // e
        64'b0000000000000000110111001101110011101101110111010000000000000000, // f
		  		  // code 0110110000
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0111000000 P
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b1111111111111111111111110000000000000000000000000000000000000000, // 2 ******
        64'b0000111111110000000011111111000000000000000000000000000000000000, // 3  **  **
        64'b0000111111110000000011111111000000000000000000000000000000000000, // 4  **  **
        64'b0000111111110000000011111111000000000000000000000000000000000000, // 5  **  **
        64'b0000111111111111111111110000000000000000000000000000000000000000, // 6  *****
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 7  **
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 8  **
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 9  **
        64'b0000111111110000000000000000000000000000000000000000000000000000, // a  **
        64'b1111111111111111000000000000000000000000000000000000000000000000, // b ****
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code 0111010000 L
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 0000
        64'b0000000000000000000000000000000000000000000000000000000000000000, // 1111
        64'b1111111111111111000000000000000000000000000000000000000000000000, // 2 ****
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 3  **
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 4  **
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 5  **
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 6  **
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 7  **
        64'b0000111111110000000000000000000000000000000000000000000000000000, // 8  **
        64'b0000111111110000000000001111000000000000000000000000000000000000, // 9  **   *
        64'b0000111111110000000011111111000000000000000000000000000000000000, // a  **  **
        64'b1111111111111111111111111111000000000000000000000000000000000000, // b *******
        64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
		  		  // code x05 placeholder
		  64'b0000000000000000010001000100010000000000000000000000000000000000, // 0
        64'b0000000000000100100010001000100001000000000000000000000000000000, // 1
        64'b0000000001001000100010000100010000000000000000000000000000000000, // 2
        64'b0000000001001010100010101010101001000000000000000000000000000000, // 3
        64'b0000010010101010101010100100101010100100000001000100010001000000, // 4
        64'b0000010001000101101010100100101010101010010010101010101001000000, // 5
        64'b0100100110011001010110100100101010101010101010101010101010100100, // 6
        64'b0000010001000101010110101010101010101010101010101010100100000000, // 7
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 8
        64'b0100010110101010101010101010101010101010101010101010010101000000, // 9
        64'b0100010110101010101010101010101010101010101010101010010101000000, // a
        64'b0000010001011010101010101010101001000101101010101010101001000000, // b
        64'b0100100101000101010101010100100101000101010110101010010000000000, // c
        64'b0100010010010100010001000100010010010100010001000100000000000000, // d
        64'b0000000000000000000000000000000000000000000000000000000000000000, // e
        64'b0000000000000000000000000000000000000000000000000000000000000000, // f
        };

	assign data = ROM[addr];

endmodule  