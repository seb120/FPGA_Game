library verilog;
use verilog.vl_types.all;
entity usb_system_mm_interconnect_0 is
    port(
        clk_clk_clk     : in     vl_logic;
        clocks_c0_clk   : in     vl_logic;
        cpu_reset_n_reset_bridge_in_reset_reset: in     vl_logic;
        sdram_reset_reset_bridge_in_reset_reset: in     vl_logic;
        cpu_data_master_address: in     vl_logic_vector(28 downto 0);
        cpu_data_master_waitrequest: out    vl_logic;
        cpu_data_master_byteenable: in     vl_logic_vector(3 downto 0);
        cpu_data_master_read: in     vl_logic;
        cpu_data_master_readdata: out    vl_logic_vector(31 downto 0);
        cpu_data_master_write: in     vl_logic;
        cpu_data_master_writedata: in     vl_logic_vector(31 downto 0);
        cpu_data_master_debugaccess: in     vl_logic;
        cpu_instruction_master_address: in     vl_logic_vector(28 downto 0);
        cpu_instruction_master_waitrequest: out    vl_logic;
        cpu_instruction_master_read: in     vl_logic;
        cpu_instruction_master_readdata: out    vl_logic_vector(31 downto 0);
        clock_crossing_io_s0_address: out    vl_logic_vector(21 downto 0);
        clock_crossing_io_s0_write: out    vl_logic;
        clock_crossing_io_s0_read: out    vl_logic;
        clock_crossing_io_s0_readdata: in     vl_logic_vector(31 downto 0);
        clock_crossing_io_s0_writedata: out    vl_logic_vector(31 downto 0);
        clock_crossing_io_s0_burstcount: out    vl_logic_vector(0 downto 0);
        clock_crossing_io_s0_byteenable: out    vl_logic_vector(3 downto 0);
        clock_crossing_io_s0_readdatavalid: in     vl_logic;
        clock_crossing_io_s0_waitrequest: in     vl_logic;
        clock_crossing_io_s0_debugaccess: out    vl_logic;
        clocks_pll_slave_address: out    vl_logic_vector(1 downto 0);
        clocks_pll_slave_write: out    vl_logic;
        clocks_pll_slave_read: out    vl_logic;
        clocks_pll_slave_readdata: in     vl_logic_vector(31 downto 0);
        clocks_pll_slave_writedata: out    vl_logic_vector(31 downto 0);
        cpu_jtag_debug_module_address: out    vl_logic_vector(8 downto 0);
        cpu_jtag_debug_module_write: out    vl_logic;
        cpu_jtag_debug_module_read: out    vl_logic;
        cpu_jtag_debug_module_readdata: in     vl_logic_vector(31 downto 0);
        cpu_jtag_debug_module_writedata: out    vl_logic_vector(31 downto 0);
        cpu_jtag_debug_module_byteenable: out    vl_logic_vector(3 downto 0);
        cpu_jtag_debug_module_waitrequest: in     vl_logic;
        cpu_jtag_debug_module_debugaccess: out    vl_logic;
        jtag_uart_avalon_jtag_slave_address: out    vl_logic_vector(0 downto 0);
        jtag_uart_avalon_jtag_slave_write: out    vl_logic;
        jtag_uart_avalon_jtag_slave_read: out    vl_logic;
        jtag_uart_avalon_jtag_slave_readdata: in     vl_logic_vector(31 downto 0);
        jtag_uart_avalon_jtag_slave_writedata: out    vl_logic_vector(31 downto 0);
        jtag_uart_avalon_jtag_slave_waitrequest: in     vl_logic;
        jtag_uart_avalon_jtag_slave_chipselect: out    vl_logic;
        keycode_s1_address: out    vl_logic_vector(1 downto 0);
        keycode_s1_write: out    vl_logic;
        keycode_s1_readdata: in     vl_logic_vector(31 downto 0);
        keycode_s1_writedata: out    vl_logic_vector(31 downto 0);
        keycode_s1_chipselect: out    vl_logic;
        sdram_s1_address: out    vl_logic_vector(24 downto 0);
        sdram_s1_write  : out    vl_logic;
        sdram_s1_read   : out    vl_logic;
        sdram_s1_readdata: in     vl_logic_vector(31 downto 0);
        sdram_s1_writedata: out    vl_logic_vector(31 downto 0);
        sdram_s1_byteenable: out    vl_logic_vector(3 downto 0);
        sdram_s1_readdatavalid: in     vl_logic;
        sdram_s1_waitrequest: in     vl_logic;
        sdram_s1_chipselect: out    vl_logic
    );
end usb_system_mm_interconnect_0;
